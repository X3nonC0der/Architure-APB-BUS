library verilog;
use verilog.vl_types.all;
entity APB_MAIN_TB is
end APB_MAIN_TB;
