library verilog;
use verilog.vl_types.all;
entity APB_slave2_TB is
end APB_slave2_TB;
